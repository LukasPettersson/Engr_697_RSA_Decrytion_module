`define DATA_WIDTH 64 //used
`define ADDR_WIDTH 6
`define TOTAL_ADDR (2 ** `ADDR_WIDTH) //used. 32
`define DATA_LENGTH 4096


module MonPro_tb();


reg clk,reset, startInput, getResults;
reg [3:0] state;
reg [4:0] exp_state;
wire [`DATA_WIDTH - 1: 0] res_out;
reg [`DATA_WIDTH - 1 : 0] m_input, e_input, n_input;
MonPro mp(.clk(clk),
          .reset(),
          .startInput(startInput),
          .getResult(),
          .m_input(m_input), //cipher text
          .e_input(e_input), // private key
          .n_input(n_input), // n
          .state(),
          .exp_state(),
          .res_out(res_out));

/* original message
1001111010011110001100111010000111100001110001010111111001011011000111010111100101100000001011111100010001011010111010100011110101111000010110001010001000010111010100101111010000110101101111111101110011100001110101001110011001101110000011011101110100011111001000010100100000011110110110101110101100001110111011011001000001111101000110000110110011000001000101011000001111000100100001010010000111101010010111100001101000011011101000110011000110110100111000100010010001001100011101011111100111011011110110101111001111111011111100000101101111101101100100010110011100011100101101111000101001100010011011011110111101100011001000110101100100100010100001111010001000000011010010010110011111001011111101110111010011000110011000111011011011000100100010010101011100110110001001001111000011001100000000010101100001001001101001010101010010000000100000110101000101101011000001000110001110111110101011010001001011100011011111101111000000010110011111101010100010011110111111110011111001111000111010110000011010001010110100100001100111101100
*/

/* encrypted message

*/
always
  #50 clk = ~clk;


initial
begin
  clk = 0;
  #50
  startInput = 1;
  #100
n_input = 64'hEAA06C6A1B82DFBB;
m_input = 64'h5B32DD707D25FCB0;
e_input = 64'h6E74641191D3CDF1;
#100
n_input = 64'h9DBCDF39485144D5;
m_input = 64'hEB961218698CF89E;
e_input = 64'h24E30DAB0E02CC43;
#100
n_input = 64'h2AA84A58A0E1708F;
m_input = 64'h1F31E0A0F55FA975;
e_input = 64'h98E325A1676F5661;
#100
n_input = 64'hBEC76F3B194537FA;
m_input = 64'hBF68A172A214EB07;
e_input = 64'hB1F84CB81B826D78;
#100
n_input = 64'h1EEBBF94EDC15519;
m_input = 64'hE99E8ECD6968F483;
e_input = 64'h1A2792E533D1502F;
#100
n_input = 64'h107E0B5CB0A1D6F8;
m_input = 64'h89F217011A7DA8B5;
e_input = 64'h63B39623CB990C60;
#100
n_input = 64'h918705100BBFD50C;
m_input = 64'h2A7E6DA76D337265;
e_input = 64'hB2412AB80208778D;
#100
n_input = 64'h923CB920D5098490;
m_input = 64'h7B9194994CA11557;
e_input = 64'hA10C5A7F76A6A346;
#100
n_input = 64'h6070683D526BC68D;
m_input = 64'hD34D7046900A8714;
e_input = 64'h73FBB168984596B0;
#100
n_input = 64'h85F91AA3CF9FA006;
m_input = 64'h292E2C056DE249AE;
e_input = 64'hEE6B160D8FF57649;
#100
n_input = 64'h8F80B52365725D12;
m_input = 64'h7E98A4A428B2F24E;
e_input = 64'h71E735F08494363B;
#100
n_input = 64'hF81A6B21B53985FF;
m_input = 64'h5A14921554696BF2;
e_input = 64'h40AF84297BBF1E91;
#100
n_input = 64'hE0BCE97AF59B468B;
m_input = 64'hBF673552129BB8FE;
e_input = 64'h9CAC839E2D957459;
#100
n_input = 64'h959ACF90FEE50B2C;
m_input = 64'h9FA29B9A365DEB1F;
e_input = 64'h81E075FA530CB570;
#100
n_input = 64'h08220E61AF5A7C08;
m_input = 64'h19EA4B4243CD9E34;
e_input = 64'hD11089654EC3FC43;
#100
n_input = 64'h8732E5420AE6D414;
m_input = 64'h254A8D1A449EBD11;
e_input = 64'h0B738D2595E4CD4B;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100
n_input = 64'h0000000000000000;
m_input = 64'h0000000000000000;
e_input = 64'h0000000000000000;
#100;
end

endmodule
