`define DATA_WIDTH 64 //used
`define ADDR_WIDTH 6
`define TOTAL_ADDR (2 ** `ADDR_WIDTH) //used. 32
`define DATA_LENGTH 4096
`define T_DATA (`DATA_LENGTH * 2) // 4096 * 2 = 8192

module constant_r_t_new_tb();

reg clk, start;
reg [`DATA_LENGTH - 1: 0] M_r;
wire [`DATA_LENGTH - 1 : 0] R_r;
wire [`DATA_LENGTH - 1 : 0] R_t;
wire done;



always #25 clk = ~clk;


initial begin
	clk = 0;
	//M_r = 1024'b0110000100010001100100000011101101011111011010110110100110111110000011000011001000011101011111010010010100111111100100011110000101001101110100000001111000001110101101101111111010001011001000001110111011100011000001001101100111101110011000110000100010100110110111000001100010101101001000001010001111000110110011001001010110110010010000100000011001111111010011111011101000011001110111101011111010100100100100110001010000000000111100101100000001111110011000000111010101100110000001000110000111011110111000101101110111000001010100100110100101110011100110100111011000011110010000010110100110101111110111011000000001010010000011110100001111011001100110000010101101000100111000001000111001001110111000110100111011100010011111010101001101111100000101110110110010110101010101100000110110000001010101110000010111000011111100111001011000000110011111000011101110001100001010110100011111101110000101100110000000010001011010101001011111000000111101110011010110101001100110101100110010011111100111111010000000111101011101101001110011111001; //Divisor
	M_r = 4096'h84c5b4763fe31d0347fc816ac16e2284c10faa4003ba33db73f7ba8e0445d656de3a5db5154ed51212093d26ac512b01f18dd1eed77c96c0084f3dd6415af341ee52bdb6d1020a15d9ed17e3cc0e95ee8d103ed3cc667e971773308cdc6b13ab2e47dc0e959f3a518cfe5cd12d5db79ba2a7ae1f3ac7652ccdf8440407295e4299901c0475491bc354c56c9a9cc9af4ec9546b439f9d01298a449ebe89d9bf020067dba8589890086a17b9af5b569643d037cdff7c240d4969d495dd81355c53f0e642f43328ad088ded3c9691eb79fa5d5f576cdeb8fc4c7b297d0b0e5e18baf320cd576d14475b349aae908fb5262cc703806984c8199921167d8fcf23cae883333218bd91a1b7f03edca7e2dcaa37f463b337d20b5d59db610487c89da11b62397bc701762741bab9f87ff50592859be3cecb8c497c68a8c24d4244ef7febe8e5b4617589a82b5a702cfa93ea5c4ed8f33418f3d4e7115804f92283868a29678a5aa33b6fe5078c5fe8f8dc3bf364eb8ac8ce8a245e6b33138131c541013d0326324dfb695ffb3a1890c78092b4d42b28fef02b9c014ea5ac06d864c2f2e39403560d97dae38d9d643c25fbb230bbd92a4aa2b410d93c4efbc8d60b21fbac78255d6807923986bb968a437d5c8dfc5eda92d864ac5db9d707107e855c384429e821a4c74803e31ba1621582283d15a9ec0806705fca161622bd795fec898f;
	#50
	start = 1;
	#50
	start = 0;
end




constant_r_t_new dut(
	.clk(clk),
	.M_r(M_r), // M is divisor
	.start(start),
	.R_r(R_r), //Remainder
	.R_t(R_t), //Remainder
	.done(done)
	);

endmodule
