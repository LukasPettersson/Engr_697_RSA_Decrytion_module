`define DATA_WIDTH 64 //used
`define ADDR_WIDTH 6
`define TOTAL_ADDR (2 ** `ADDR_WIDTH) //used. 32
`define DATA_LENGTH 4096


module MonPro_tb();


reg clk,reset, startInput, getResults;
reg [3:0] state;
reg [4:0] exp_state;
wire [`DATA_WIDTH - 1: 0] res_out;
reg [`DATA_WIDTH - 1 : 0] m_input, e_input, n_input;
MonPro mp(.clk(clk),
          .reset(),
          .startInput(startInput),
          .getResult(),
          .m_input(m_input), //cipher text
          .e_input(e_input), // private key
          .n_input(n_input), // n
          .state(),
          .exp_state(),
          .res_out(res_out));

/* original message
1001111010011110001100111010000111100001110001010111111001011011000111010111100101100000001011111100010001011010111010100011110101111000010110001010001000010111010100101111010000110101101111111101110011100001110101001110011001101110000011011101110100011111001000010100100000011110110110101110101100001110111011011001000001111101000110000110110011000001000101011000001111000100100001010010000111101010010111100001101000011011101000110011000110110100111000100010010001001100011101011111100111011011110110101111001111111011111100000101101111101101100100010110011100011100101101111000101001100010011011011110111101100011001000110101100100100010100001111010001000000011010010010110011111001011111101110111010011000110011000111011011011000100100010010101011100110110001001001111000011001100000000010101100001001001101001010101010010000000100000110101000101101011000001000110001110111110101011010001001011100011011111101111000000010110011111101010100010011110111111110011111001111000111010110000011010001010110100100001100111101100
*/

/* encrypted message

*/
always
  #50 clk = ~clk;


initial
begin
  clk = 0;
  #50
  startInput = 1;
  #100
n_input = 64'hE29A87C176A78B35;
m_input = 64'h384CB8DCF02466CE;
e_input = 64'h1A32639C11288001;
#100
n_input = 64'h96DC65A491BFACCF;
m_input = 64'hAFE16C009C180116;
e_input = 64'h55A83A5C8979F547;
#100
n_input = 64'h912B843C829D66CD;
m_input = 64'h7CF0F85F8D0E3DBB;
e_input = 64'hAFE6DEF43224F223;
#100
n_input = 64'h6A9B8743E2AC3B9E;
m_input = 64'h047FA9F23C85C959;
e_input = 64'h2B01B3BF40A7B474;
#100
n_input = 64'hCB623CDB9994BD5F;
m_input = 64'hB2A22C3B49EA3C8C;
e_input = 64'h71066FE1504B6DCF;
#100
n_input = 64'h6104CCF491C408C7;
m_input = 64'h3B84DBFF6642915A;
e_input = 64'h82BE1C4144528D50;
#100
n_input = 64'h77503DA8686D4D67;
m_input = 64'h931B325D4F2C2F83;
e_input = 64'hBF5A874406653F01;
#100
n_input = 64'h3C2F2CC478B9A4EA;
m_input = 64'h825D6EDF1FB3960C;
e_input = 64'h2D94C1AD4D63009B;
#100
n_input = 64'h9863A2A0DD158527;
m_input = 64'hA8BF244C51618B96;
e_input = 64'h5B32A1235B4FA3B8;
#100
n_input = 64'h88857AE67E466429;
m_input = 64'h9A13B4F8B7C088AA;
e_input = 64'h1BD907DB8069D369;
#100
n_input = 64'hF50EED41AB792974;
m_input = 64'h9CD81AEAE5CC806E;
e_input = 64'hED2B316514075437;
#100
n_input = 64'h89ADFF6ED1E584EE;
m_input = 64'hCE66E06A4EFA53B2;
e_input = 64'hC51DD6ED3797DA73;
#100
n_input = 64'h9E45B3A5B3EBBD09;
m_input = 64'h6AE92E9318452B0A;
e_input = 64'h69C65B26108411F7;
#100
n_input = 64'h068D5609ABCCD6A0;
m_input = 64'h55BE19DB7149BDE6;
e_input = 64'hE9961FA1CCE712CD;
#100
n_input = 64'hB637CC375EA40B10;
m_input = 64'h1A607A5829B8986C;
e_input = 64'hCD7CDEB546BB8BDC;
#100
n_input = 64'h5FB8536C1E49899B;
m_input = 64'h7FEBC9BA3017691E;
e_input = 64'h0D1CDB25A563A9B1;
#100
n_input = 64'h5D908F8EB8C215B0;
m_input = 64'h1829C1D58338BA25;
e_input = 64'h77C3CC50BC06C60E;
#100
n_input = 64'hFC3354F4739A0DFE;
m_input = 64'h175B16D02F9FF61A;
e_input = 64'h2E6E4769CF3E3B43;
#100
n_input = 64'h24BCE3AF4132A935;
m_input = 64'hEB069047E4D87265;
e_input = 64'h287CD1973745D4C3;
#100
n_input = 64'h06DA7B7639C96814;
m_input = 64'h3DC5FF45640D8A14;
e_input = 64'h716E6F60345D608A;
#100
n_input = 64'h759198AB32136F4F;
m_input = 64'hF8A01A7B38989CAB;
e_input = 64'h72A400954AA6B702;
#100
n_input = 64'h20E1D5B87C751B1C;
m_input = 64'h35E26587325563EA;
e_input = 64'h6AB6F267D6B02477;
#100
n_input = 64'hC887ABFB984B4A08;
m_input = 64'hFD1DDA2BF6F37690;
e_input = 64'hB8276FBBC3B49E8F;
#100
n_input = 64'h109EFB4AFFA904F3;
m_input = 64'h9CFF957BA0FE423C;
e_input = 64'h25D6097321BFE47B;
#100
n_input = 64'h07892FB0E121F76D;
m_input = 64'h8113C31851909ACE;
e_input = 64'h954D5CBE9344C91A;
#100
n_input = 64'h1C7D7C40ABC74199;
m_input = 64'h8031796DEB142868;
e_input = 64'hBB4A13B45E18112C;
#100
n_input = 64'h3CFBD9DD0F63B0CE;
m_input = 64'hD18943458FF58E69;
e_input = 64'h2D39CABAE504CA87;
#100
n_input = 64'h4FDFB937D870D834;
m_input = 64'hBA7AE23C8CF1F971;
e_input = 64'h3C6533377B5A17EB;
#100
n_input = 64'h0D74E1B07D44A9F9;
m_input = 64'hF7A23F8618A388C4;
e_input = 64'hD0903684585A7391;
#100
n_input = 64'h2E6EE2C622CBB96D;
m_input = 64'h4559367361B0477C;
e_input = 64'h2F849AB4355AEC72;
#100
n_input = 64'h952A54C69107E72F;
m_input = 64'hF8243598DB6A1AAA;
e_input = 64'h7688945F69521137;
#100
n_input = 64'hCF13F2B8A92D537D;
m_input = 64'h457D5136284FA11F;
e_input = 64'h099FA0FCC75B62B1;
#100
n_input = 64'h6CB07B526BB8EE0A;
m_input = 64'hA389AF082C4A920E;
e_input = 64'hF2138E05DE0C4C4D;
#100
n_input = 64'h60A5A53A845713AA;
m_input = 64'h471DFC34E3B60DF8;
e_input = 64'hF880C33389083C37;
#100
n_input = 64'h007A60D976E815EC;
m_input = 64'h19971A0D19995E55;
e_input = 64'h9D48755952FD2206;
#100
n_input = 64'h4440EFAE4CD23653;
m_input = 64'hFEF3744A351C0AB0;
e_input = 64'hAF4C2A303243E815;
#100
n_input = 64'h58AC05202E0D820C;
m_input = 64'h4A07D7EADF490DAE;
e_input = 64'hC94338D31E8564E6;
#100
n_input = 64'h6261F9EEFCC831CE;
m_input = 64'hF4F5F997EBBEAE45;
e_input = 64'h82D949ADE52591FB;
#100
n_input = 64'h4CFC58F4ACDC83C9;
m_input = 64'h97AB88545360A058;
e_input = 64'hE07627ABC4B9F7E1;
#100
n_input = 64'h7122BA2BF761418B;
m_input = 64'h0995F5864DAF1FA4;
e_input = 64'h642270B1308BD385;
#100
n_input = 64'h48B18D07BE889015;
m_input = 64'h77E1B66DCA39B574;
e_input = 64'h3F333D5D24379B87;
#100
n_input = 64'h0795E139C4E4C558;
m_input = 64'h0417478986835888;
e_input = 64'h9DFBAA601865778B;
#100
n_input = 64'h1986BD1C574498F9;
m_input = 64'hFDF31C39EF896A8A;
e_input = 64'h37745B976992A8BC;
#100
n_input = 64'hE7CF05CF53E4B975;
m_input = 64'hD3836936D7D2F70C;
e_input = 64'hDD79FB70E2B39A2E;
#100
n_input = 64'hB6B924C1FB22470F;
m_input = 64'h3358687AEE7ABE9E;
e_input = 64'h0015FB8C06BDE91A;
#100
n_input = 64'hE96DD6A8A42F58D0;
m_input = 64'h0E187F8D8E77E207;
e_input = 64'hA312B799FE729F0A;
#100
n_input = 64'hB1467B400D6964A1;
m_input = 64'h4EDB2627F24DE9AC;
e_input = 64'hA4D1E6B3B48139EE;
#100
n_input = 64'h026B4C6F739DC0C3;
m_input = 64'h8012A39267059AA3;
e_input = 64'h59B12A4EEA151FE6;
#100
n_input = 64'h4913159E219826CF;
m_input = 64'hCE5AB278157B85A7;
e_input = 64'h89B873245C0B0FC8;
#100
n_input = 64'h2D28A12AF9F18CED;
m_input = 64'h098E6109F340201D;
e_input = 64'hD8AD4716B04F95B5;
#100
n_input = 64'h471FF21A5C962577;
m_input = 64'hADE2DFD13CCA2165;
e_input = 64'h8E7E0B582839432B;
#100
n_input = 64'h703E900A0FEB6A62;
m_input = 64'h9C5F886A8433CE32;
e_input = 64'hE5B8D9354EDCCEE1;
#100
n_input = 64'hE7BAD3BCFC602DE2;
m_input = 64'h0164DACF766F390B;
e_input = 64'h9779A98AEAA04A25;
#100
n_input = 64'h9D93EF6A83E3D697;
m_input = 64'h0CD923D9419C9DDA;
e_input = 64'h20B5C7D3BCD6FF82;
#100
n_input = 64'h32F42A6E479EC1EB;
m_input = 64'hAC6268155331E97F;
e_input = 64'h68BEF82700968ED1;
#100
n_input = 64'hC2633ED13AAEDB6D;
m_input = 64'hA6253EA4154598DB;
e_input = 64'h965B0069AADCA845;
#100
n_input = 64'h4A112D3CEB858232;
m_input = 64'h0FF4658A78F00EBF;
e_input = 64'hC34357CA6A34DED7;
#100
n_input = 64'hD0476589DB421C4B;
m_input = 64'h6F881268A082A973;
e_input = 64'h9FF8213E6D6B4DFA;
#100
n_input = 64'h9641EC994548E33E;
m_input = 64'hA0BFC53942108E36;
e_input = 64'hE6B79A630556244B;
#100
n_input = 64'hD233E515FC3DB05D;
m_input = 64'hE2322833429EC4D1;
e_input = 64'h0C1D44C6FC138BAD;
#100
n_input = 64'h94A5D1192F1E2463;
m_input = 64'hE2CF2F80C158D2C7;
e_input = 64'hC1166548A001E55E;
#100
n_input = 64'h695490240ECE5D0F;
m_input = 64'h5A6C78A3F83151EA;
e_input = 64'hDEA9BAC37D01561B;
#100
n_input = 64'h5F0E520DFF1EA7DF;
m_input = 64'h781B85403EFD11B6;
e_input = 64'hE32286CBA9D87379;
#100
n_input = 64'h5FAF79A3517B1A13;
m_input = 64'h0DAB8BDAFE504EEB;
e_input = 64'h28B6D3BD287886F9;
#100;
end

endmodule
