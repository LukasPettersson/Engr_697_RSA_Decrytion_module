module n0prime_new_tb();



reg [2047:0] p,q;
wire [2047:0] t,qinv;
reg start, clk;
wire done;

  n0prime dut(
              .p(p),
              .q(q),
              .t(t),
              .qinv(qinv),
              .start(start),
              .clk(clk),
              .done(done));

  always
    #5 clk = ~clk;


  initial begin
    clk <=0;
    //p has to be smaller than q to get the right answer
    //n = 110620781787982559320879672277187232847059370855697531032471456562776629662302244635541635743974443111884235645205863300149086076806673694355442778484112581750287392626037519520354184007761932200792383173427168395884973735814267160431334221012878580946600314337283120169876076782148446769399989029866652585707
    q <= 2048'd110620781787982559320879672277187232847059370855697531032471456562776629662302244635541635743974443111884235645205863300149086076806673694355442778484112581750287392626037519520354184007761932200792383173427168395884973735814267160431334221012878580946600314337283120169876076782148446769399989029866652585707;
    p <= 2048'd4294967296;
    start <= 1;
    #10
    start <= 0;
  end


endmodule
