`define DATA_WIDTH 32 //used
`define ADDR_WIDTH 5
`define TOTAL_ADDR (2 ** `ADDR_WIDTH) //used. 32
`define DATA_LENGTH 1024


module MonPro_tb();


reg clk,reset, startInput, getResults;
reg [3:0] state;
reg [4:0] exp_state;
wire [31 : 0] res_out;
reg [`DATA_WIDTH - 1 : 0] m_input, e_input, n_input;
MonPro mp(.clk(clk),
          .reset(),
          .startInput(startInput),
          .getResult(),
          .m_input(m_input), //cipher text
          .e_input(e_input), // private key
          .n_input(n_input), // n
          .state(),
          .exp_state(),
          .res_out(res_out));

/* original message
1001111010011110001100111010000111100001110001010111111001011011000111010111100101100000001011111100010001011010111010100011110101111000010110001010001000010111010100101111010000110101101111111101110011100001110101001110011001101110000011011101110100011111001000010100100000011110110110101110101100001110111011011001000001111101000110000110110011000001000101011000001111000100100001010010000111101010010111100001101000011011101000110011000110110100111000100010010001001100011101011111100111011011110110101111001111111011111100000101101111101101100100010110011100011100101101111000101001100010011011011110111101100011001000110101100100100010100001111010001000000011010010010110011111001011111101110111010011000110011000111011011011000100100010010101011100110110001001001111000011001100000000010101100001001001101001010101010010000000100000110101000101101011000001000110001110111110101011010001001011100011011111101111000000010110011111101010100010011110111111110011111001111000111010110000011010001010110100100001100111101100
*/

/* encrypted message

*/
always
  #50 clk = ~clk;


initial
begin
  clk = 0;
  #50
  startInput = 1;
  #100
  n_input = 32'h8B9496E5;
m_input = 32'h00000005;
e_input = 32'h00010001;
#100
n_input = 32'h5F06287C;
m_input = 32'h00000000;
e_input = 32'h00000000;
#100
n_input = 32'h31988514;
m_input = 32'h00000000;
e_input = 32'h00000000;
#100
n_input = 32'hF96F9A0B;
m_input = 32'h00000000;
e_input = 32'h00000000;
#100
n_input = 32'h098EC99C;
m_input = 32'h00000000;
e_input = 32'h00000000;
#100
n_input = 32'hCE60DEFE;
m_input = 32'h00000000;
e_input = 32'h00000000;
#100
n_input = 32'h7B044519;
m_input = 32'h00000000;
e_input = 32'h00000000;
#100
n_input = 32'h197CBC98;
m_input = 32'h00000000;
e_input = 32'h00000000;
#100
n_input = 32'h8C547944;
m_input = 32'h00000000;
e_input = 32'h00000000;
#100
n_input = 32'h528B17F6;
m_input = 32'h00000000;
e_input = 32'h00000000;
#100
n_input = 32'h024D981B;
m_input = 32'h00000000;
e_input = 32'h00000000;
#100
n_input = 32'h9397F02E;
m_input = 32'h00000000;
e_input = 32'h00000000;
#100
n_input = 32'h13F7DBF4;
m_input = 32'h00000000;
e_input = 32'h00000000;
#100
n_input = 32'h65D03E3B;
m_input = 32'h00000000;
e_input = 32'h00000000;
#100
n_input = 32'hE3DA97CB;
m_input = 32'h00000000;
e_input = 32'h00000000;
#100
n_input = 32'hE728F169;
m_input = 32'h00000000;
e_input = 32'h00000000;
#100
n_input = 32'hA0FA5221;
m_input = 32'h00000000;
e_input = 32'h00000000;
#100
n_input = 32'h6FB2A652;
m_input = 32'h00000000;
e_input = 32'h00000000;
#100
n_input = 32'h4F8EA1A0;
m_input = 32'h00000000;
e_input = 32'h00000000;
#100
n_input = 32'h5ABE53AE;
m_input = 32'h00000000;
e_input = 32'h00000000;
#100
n_input = 32'h12A3EAD3;
m_input = 32'h00000000;
e_input = 32'h00000000;
#100
n_input = 32'h8C4CB074;
m_input = 32'h00000000;
e_input = 32'h00000000;
#100
n_input = 32'h1487CE4E;
m_input = 32'h00000000;
e_input = 32'h00000000;
#100
n_input = 32'h5BC6D48D;
m_input = 32'h00000000;
e_input = 32'h00000000;
#100
n_input = 32'h2F604851;
m_input = 32'h00000000;
e_input = 32'h00000000;
#100
n_input = 32'h2C34DF98;
m_input = 32'h00000000;
e_input = 32'h00000000;
#100
n_input = 32'h0AD14479;
m_input = 32'h00000000;
e_input = 32'h00000000;
#100
n_input = 32'hC1526B25;
m_input = 32'h00000000;
e_input = 32'h00000000;
#100
n_input = 32'h0357F18C;
m_input = 32'h00000000;
e_input = 32'h00000000;
#100
n_input = 32'hD18C0F37;
m_input = 32'h00000000;
e_input = 32'h00000000;
#100
n_input = 32'hA346920B;
m_input = 32'h00000000;
e_input = 32'h00000000;
#100
n_input = 32'hA938A368;
m_input = 32'h00000000;
e_input = 32'h00000000;
#100; 
end

endmodule
