`define DATA_WIDTH 64 //used
`define ADDR_WIDTH 6
`define TOTAL_ADDR (2 ** `ADDR_WIDTH) //used. 32
`define DATA_LENGTH 4096


module MonPro_tb();


reg clk,reset, startInput, getResults;
reg [3:0] state;
reg [4:0] exp_state;
wire [`DATA_WIDTH - 1: 0] res_out;
reg [`DATA_WIDTH - 1 : 0] m_input, e_input, n_input;
MonPro mp(.clk(clk),
          .reset(),
          .startInput(startInput),
          .getResult(),
          .m_input(m_input), //cipher text
          .e_input(e_input), // private key
          .n_input(n_input), // n
          .state(),
          .exp_state(),
          .res_out(res_out));

/* original message
1001111010011110001100111010000111100001110001010111111001011011000111010111100101100000001011111100010001011010111010100011110101111000010110001010001000010111010100101111010000110101101111111101110011100001110101001110011001101110000011011101110100011111001000010100100000011110110110101110101100001110111011011001000001111101000110000110110011000001000101011000001111000100100001010010000111101010010111100001101000011011101000110011000110110100111000100010010001001100011101011111100111011011110110101111001111111011111100000101101111101101100100010110011100011100101101111000101001100010011011011110111101100011001000110101100100100010100001111010001000000011010010010110011111001011111101110111010011000110011000111011011011000100100010010101011100110110001001001111000011001100000000010101100001001001101001010101010010000000100000110101000101101011000001000110001110111110101011010001001011100011011111101111000000010110011111101010100010011110111111110011111001111000111010110000011010001010110100100001100111101100
*/

/* encrypted message

*/
always
  #50 clk = ~clk;


initial
begin
  clk = 0;
  #50
  startInput = 1;
  #100
  n_input = 64'h31986649780FA7EF;
  m_input = 64'h66FFE53674D8AD58;
  e_input = 64'h53CE65B0C1F8D001;
  #100
  n_input = 64'hF72D58F492D5B712;
  m_input = 64'hEADAC2DE0A05C170;
  e_input = 64'hEFE9341764279FE5;
  #100
  n_input = 64'h18253BC33F3BE25A;
  m_input = 64'h1B171B253F0BEA91;
  e_input = 64'hB913C495911B3CC9;
  #100
  n_input = 64'hC292E93436516642;
  m_input = 64'h1E1FA15837734C85;
  e_input = 64'hA958846B3CC64120;
  #100
  n_input = 64'h6B6CD6F10C0573BF;
  m_input = 64'h457F720E4793E2D3;
  e_input = 64'h8E26A0F54BB32144;
  #100
  n_input = 64'h2641CA9F9C3B9693;
  m_input = 64'hC2871421D713373F;
  e_input = 64'h43A638947FC665E8;
  #100
  n_input = 64'hC181EB3B2B021B2C;
  m_input = 64'hA86F9FACFDB73506;
  e_input = 64'h82CF2A5147E67461;
  #100
  n_input = 64'h833016EACFF2E19D;
  m_input = 64'hF64F2B50C4F5532C;
  e_input = 64'hC859DB3DFF4891E7;
  #100
  n_input = 64'hC93C2EE0FF66536B;
  m_input = 64'h6AE29859C802A04E;
  e_input = 64'h0645BE41DA3F9908;
  #100
  n_input = 64'h842317807D7011DE;
  m_input = 64'h7E88A2D1583ED3B7;
  e_input = 64'h3ABF521F963EF914;
  #100
  n_input = 64'hC35FB76C946A4EB3;
  m_input = 64'hCBDF5825F60B4E26;
  e_input = 64'hA5F78E5D50662666;
  #100
  n_input = 64'h4B472BCC22831A71;
  m_input = 64'h7F0540B03487460D;
  e_input = 64'hB621101DECCF9330;
  #100
  n_input = 64'hEB94791004DD4A01;
  m_input = 64'hEAA8D90F21201DED;
  e_input = 64'h863AAA5075AF937D;
  #100
  n_input = 64'hB04F0848CCF5D6DF;
  m_input = 64'h98B55DE719A0C474;
  e_input = 64'h26D20AFED0081B77;
  #100
  n_input = 64'h5CC5B1A92CDC6FB9;
  m_input = 64'h7613510835A6C1FE;
  e_input = 64'h9B3C8C763763381E;
  #100
  n_input = 64'hCED8117AA872DD99;
  m_input = 64'h1269B27176B50B29;
  e_input = 64'hA32570D9D8F5B827;
  #100
  n_input = 64'h492FB0044D92E5B8;
  m_input = 64'hCA840F37CF2CFCB0;
  e_input = 64'hA5B4B42168EC5B21;
  #100
  n_input = 64'h6C2440EAFF931B46;
  m_input = 64'h0AA4A397D65B19B4;
  e_input = 64'h984FD41258445E24;
  #100
  n_input = 64'h9848B4008D99267D;
  m_input = 64'h7C7CFB63F9A9BFEA;
  e_input = 64'hAE3096B67C38BFB9;
  #100
  n_input = 64'h2B7B87C97C50B438;
  m_input = 64'h1B90C02A28352C18;
  e_input = 64'hBD83004A80AA4CBA;
  #100
  n_input = 64'h9328867C891D2055;
  m_input = 64'h033B749A7C926BA2;
  e_input = 64'hBD6603F17C2204C4;
  #100
  n_input = 64'h9E6D8EE5DE47A215;
  m_input = 64'hC6F8EB6E107A5807;
  e_input = 64'hE781B63E36302B73;
  #100
  n_input = 64'hC04B8E4D9C300E8A;
  m_input = 64'h8ACC0E4220633000;
  e_input = 64'h33545844CE1A1C05;
  #100
  n_input = 64'h8FD2314AC1B7B88A;
  m_input = 64'hE3C0463F02B0D81E;
  e_input = 64'h2B7894DAB873AF92;
  #100
  n_input = 64'h510B5AB30C7A05AB;
  m_input = 64'hB9A7C3FAED3B8702;
  e_input = 64'h952B8617BE2B8572;
  #100
  n_input = 64'h3CC0696E377148CF;
  m_input = 64'hE2E55087F04432C6;
  e_input = 64'hCDAF50ECBC131004;
  #100
  n_input = 64'h73AA9022D3BC7027;
  m_input = 64'h1D040DA3029B0F0B;
  e_input = 64'h2159E5878336B5A5;
  #100
  n_input = 64'hEB1DC6B4253A8FF9;
  m_input = 64'hDDA7961799FD0ABF;
  e_input = 64'h9FEF5244958F9BAF;
  #100
  n_input = 64'h92B7365744152DE3;
  m_input = 64'h9F7673B83E22CAFD;
  e_input = 64'hFCBE2651EB1AB239;
  #100
  n_input = 64'h5DC3FB8121152C6E;
  m_input = 64'h5D5561C26CF94BC9;
  e_input = 64'hD9576C266F2D2789;
  #100
  n_input = 64'hC8B4965B44B16127;
  m_input = 64'hF99BE5226AEF0FBE;
  e_input = 64'hEB95B67426F9C805;
  #100
  n_input = 64'h71B36E4E97B2B6AA;
  m_input = 64'h56C4E621FD4673BC;
  e_input = 64'h3405B314169D5654;
  #100
  n_input = 64'h3773E72DFAF51A44;
  m_input = 64'h2938E1AB4345EA2D;
  e_input = 64'hA617145F9CA84F83;
  #100
  n_input = 64'h12C58A41D9185ED3;
  m_input = 64'h636BB2F6287372DE;
  e_input = 64'hBC86BFCC14949A0E;
  #100
  n_input = 64'hB4A1B8A107976929;
  m_input = 64'h8D2267936B93DA71;
  e_input = 64'h20DF29F3958617BF;
  #100
  n_input = 64'h3F6065BAC3BAD5BE;
  m_input = 64'hBBD3A62849868B87;
  e_input = 64'hF3F26C2014EF7A4E;
  #100
  n_input = 64'h4FD4E6B50D8771AD;
  m_input = 64'h3A8AD22E4EACC93C;
  e_input = 64'hC3FB4F9C3289E96F;
  #100
  n_input = 64'hE644EF1092578F05;
  m_input = 64'h33349143E4D4F976;
  e_input = 64'hB7B38A7800B7EA5A;
  #100
  n_input = 64'h9B1EC43750FAC855;
  m_input = 64'hB74B4F87348FBBCD;
  e_input = 64'hACD80A997FA3E50B;
  #100
  n_input = 64'h20478B3614761E14;
  m_input = 64'h0E3281D38C3FD265;
  e_input = 64'hAC64A3AE6D6C8B40;
  #100
  n_input = 64'h4DF35870F75A313F;
  m_input = 64'hE9C96ED2A228B5A2;
  e_input = 64'h19AAF071FA3F8383;
  #100
  n_input = 64'h65ACF8FF71A1C1C5;
  m_input = 64'hA5AA27AB3C9CEE8F;
  e_input = 64'hB4E0F11C1ED4B330;
  #100
  n_input = 64'hC5F703EFE6F778C1;
  m_input = 64'h86FD4D82111B60C4;
  e_input = 64'hDE330F6644E584A6;
  #100
  n_input = 64'h25E53D3489DD4133;
  m_input = 64'hA1862F148D389449;
  e_input = 64'h59DC95D044B3621E;
  #100
  n_input = 64'hC5A898EC42287D2D;
  m_input = 64'hB47EC4EF748F02EA;
  e_input = 64'h6D5AC7032F0FAF77;
  #100
  n_input = 64'hAEB26D84217DF056;
  m_input = 64'hC120B92584A1D711;
  e_input = 64'hB249BEE9C172DF39;
  #100
  n_input = 64'h40A2CE288DD6E0B6;
  m_input = 64'hE20BC5F1837B62E8;
  e_input = 64'hC34861FC89A81837;
  #100
  n_input = 64'h63BDCA84817B1CB3;
  m_input = 64'h8D0AA83BFEC6D7D7;
  e_input = 64'hA9FC38EB12FF5417;
  #100
  n_input = 64'hAF3B140EFB7B9B03;
  m_input = 64'h442868DF3A6CB5FA;
  e_input = 64'h7ED58174497D8105;
  #100
  n_input = 64'h51AE4C8852E02CC1;
  m_input = 64'hEB46C6DAF04D6EAF;
  e_input = 64'hE2A4CE987EA2F497;
  #100
  n_input = 64'h6D361217050DAF4B;
  m_input = 64'h1DD875D8D486397A;
  e_input = 64'h5016BF265F53E625;
  #100
  n_input = 64'h835553F36D581768;
  m_input = 64'h9BE32973BD001A28;
  e_input = 64'h0390A603748D61DF;
  #100
  n_input = 64'hB54A599AF098A349;
  m_input = 64'hB51D835F084C5444;
  e_input = 64'h5C5EA928CB37594F;
  #100
  n_input = 64'h8366EF211228C649;
  m_input = 64'h58AFDFB0D29355A5;
  e_input = 64'h6DAD178B703FA7D3;
  #100
  n_input = 64'hBEFA5E540AD9C2D6;
  m_input = 64'h88B59B7E2319299F;
  e_input = 64'hE6D02A6EFC1B6AC0;
  #100
  n_input = 64'h45700BEE555B9A06;
  m_input = 64'h6BE33DFAAECD58DD;
  e_input = 64'hCA6EE6F5313A6881;
  #100
  n_input = 64'h9A4468F023A878C3;
  m_input = 64'hD0710EB9BECF478B;
  e_input = 64'h06DCD1BC3254E8B8;
  #100
  n_input = 64'hE55AF53985E0AFCA;
  m_input = 64'hC6B77D331859C67D;
  e_input = 64'hB9F25E1268CDF190;
  #100
  n_input = 64'hC6355D36B57BE7AF;
  m_input = 64'hE83B349F92DBD758;
  e_input = 64'h3ECDC210CDC83914;
  #100
  n_input = 64'hF787D0D9432C12B6;
  m_input = 64'h4E4545515289F664;
  e_input = 64'hF7096FD992859E35;
  #100
  n_input = 64'hB731D363B014C408;
  m_input = 64'hB9C23FB30A33C932;
  e_input = 64'h014BB697408117CB;
  #100
  n_input = 64'hA3A2A6D7CF0A6263;
  m_input = 64'hB80AF7012DD78FE9;
  e_input = 64'hD9E7AC6B310B7B66;
  #100
  n_input = 64'h268BE6C36F0DB3B7;
  m_input = 64'h0D112F0A4886EF73;
  e_input = 64'h61C9BC5917903164;
  #100
  n_input = 64'hBE0B663C1CB96D9C;
  m_input = 64'h00039091796AE075;
  e_input = 64'h95956362ED39068D;
  #100;
end

endmodule
