module r_tb;

reg [1023:0] n;
reg clk, go;
wire [1023:0 ] ans;
wire [31:0] out;
r dut(.clk(clk), .go(go), .out(out));


always 
	#5 clk = ~clk;

	
initial begin
	clk = 0;
end

initial begin
	//n <= 1024'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	#15 go <= 1'b1;
end


endmodule
