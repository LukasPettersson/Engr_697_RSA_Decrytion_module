module MonPro_tb();


endmodule
