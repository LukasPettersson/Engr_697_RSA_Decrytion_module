module n0prime512_test;


reg [511:0] p,q;
wire [511:0] qinv, t;
reg clk,start;

 
n0prime512 dut(.q(q), .p(p), .t(t), .qinv(qinv), .clk(clk), .start(start));

/*
module n0prime(
			input  [31:0] q,p,
			output reg [31:0] qinv,
			input clk, start

*/

initial begin
	clk = 1'b1;
	start = 1'b0;
	p = 512'b0;
	q = 512'b0;
	
end

always begin
	#5 clk = ~clk;
	
end

initial
	begin
		$display("32'h0020 mod 32'h0016=%d",32'h0020 % 32'h0016);
		start = 1;
		//prime numbers (decimal)
		//p = 12889978550408541482772392516347090086328095581238914691443603501141658826038386152838464768711411078039955682544411327163774464365707463902628180515854417
		//q = 9526043210839685188726909141078919438064380825445233817716885796932211500901402250093422670036730581126527776573217006582288885625211747918571300192768553
		p = 512'hF61CE7187CC09E35C7B981BAC4051572E25699BD73E15D991B3005EA8AC0CDCB61502E139FBDE8A0D307D15A9C1EE005228B3DD9B059A2480C32D3AC5EA39851;  
		q = 512'hB5E2544C3995BD314B33973748EE1F0EF60A557B26DA2ADDB684A0C990FEE804B7D233C11959B5C633DCE5F79747613330AF6EA2CFB3C5020A1067E31887D229;  	
		
		repeat(2)@(posedge clk);
		start = 0;
		#100000


		$finish;
	 end

endmodule
