module dbs_r_tb();
	

	reg [1025:0] dividend;
	reg [1023 :0] divisor;
	reg clk;
	wire [1023:0] remainder, quotient;
	reg [12:0] num;
	wire done;
	reg start;

	dbs_r dut(.start(start), .clk(clk),.dividend(dividend),.divisor(divisor),.outputcount(quotient),.remainder(remainder),.done(done));
	
	always
		#25 clk = ~clk;
	
	initial begin
		clk = 0;
		start = 1'b1;
		num = 11'd1024;
		dividend = 1'b1 << num;
		divisor = 1024'b0110000100010001100100000011101101011111011010110110100110111110000011000011001000011101011111010010010100111111100100011110000101001101110100000001111000001110101101101111111010001011001000001110111011100011000001001101100111101110011000110000100010100110110111000001100010101101001000001010001111000110110011001001010110110010010000100000011001111111010011111011101000011001110111101011111010100100100100110001010000000000111100101100000001111110011000000111010101100110000001000110000111011110111000101101110111000001010100100110100101110011100110100111011000011110010000010110100110101111110111011000000001010010000011110100001111011001100110000010101101000100111000001000111001001110111000110100111011100010011111010101001101111100000101110110110010110101010101100000110110000001010101110000010111000011111100111001011000000110011111000011101110001100001010110100011111101110000101100110000000010001011010101001011111000000111101110011010110101001100110101100110010011111100111111010000000111101011101101001110011111001;
		
	end
	
endmodule
//0110000100010001100100000011101101011111011010110110100110111110000011000011001000011101011111010010010100111111100100011110000101001101110100000001111000001110101101101111111010001011001000001110111011100011000001001101100111101110011000110000100010100110110111000001100010101101001000001010001111000110110011001001010110110010010000100000011001111111010011111011101000011001110111101011111010100100100100110001010000000000111100101100000001111110011000000111010101100110000001000110000111011110111000101101110111000001010100100110100101110011100110100111011000011110010000010110100110101111110111011000000001010010000011110100001111011001100110000010101101000100111000001000111001001110111000110100111011100010011111010101001101111100000101110110110010110101010101100000110110000001010101110000010111000011111100111001011000000110011111000011101110001100001010110100011111101110000101100110000000010001011010101001011111000000111101110011010110101001100110101100110010011111100111111010000000111101011101101001110011111001;