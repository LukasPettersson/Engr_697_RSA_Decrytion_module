module secondaryInputTop();



/*
all:
start

n0prime:
input p, q
output t, qinv

r:
input p, q
output: 

insantiate n0prime, r, t
*/

always (@posedge clk)


endmodule
