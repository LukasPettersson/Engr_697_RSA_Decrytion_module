module shiftIn_tb;

reg clk;
reg [7:0] data;

wire [511:0] outputReg;

shiftIn dut(	.data(data), 
				.clk(clk), 
				.outputReg(outputReg)
			);

			
			
always  
	#5 clk = ~clk;

initial begin
	clk <= 0;

	
end

initial begin
		
	data <= 8'b1111111111111111;
	#15
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;

	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;

	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
	#10
	data <= 8'b1111111111111111;
end
endmodule
